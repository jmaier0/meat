
.PARAM ref='supp/2' sh='supp/2'
.PARAM opamp_amplification=-50
.PARAM R_A=10meg
.PARAM R_B=4meg
.PARAM C_0=10pF
.PARAM R_0=5
